// CPU.v

// Generated using ACDS version 13.1 162 at 2019.12.10.17:15:23

`timescale 1 ps / 1 ps
module CPU (
		input  wire       clk_clk,                                //                             clk.clk
		input  wire       reset_reset_n,                          //                           reset.reset_n
		output wire       lcd_0_conduit_end_export,               //               lcd_0_conduit_end.export
		output wire       lcd_0_conduit_end_1_export,             //             lcd_0_conduit_end_1.export
		output wire       lcd_0_conduit_end_2_export,             //             lcd_0_conduit_end_2.export
		output wire [7:0] lcd_0_conduit_end_3_export,             //             lcd_0_conduit_end_3.export
		output wire       led_external_connection_export,         //         led_external_connection.export
		input  wire       jumpbutton_external_connection_export,  //  jumpbutton_external_connection.export
		input  wire       pausebutton_external_connection_export  // pausebutton_external_connection.export
	);

	wire  [31:0] nios2_qsys_0_custom_instruction_master_result;                                   // nios2_qsys_0_custom_instruction_master_translator:ci_slave_result -> nios2_qsys_0:E_ci_result
	wire   [4:0] nios2_qsys_0_custom_instruction_master_b;                                        // nios2_qsys_0:D_ci_b -> nios2_qsys_0_custom_instruction_master_translator:ci_slave_b
	wire   [4:0] nios2_qsys_0_custom_instruction_master_c;                                        // nios2_qsys_0:D_ci_c -> nios2_qsys_0_custom_instruction_master_translator:ci_slave_c
	wire         nios2_qsys_0_custom_instruction_master_done;                                     // nios2_qsys_0_custom_instruction_master_translator:ci_slave_multi_done -> nios2_qsys_0:E_ci_multi_done
	wire         nios2_qsys_0_custom_instruction_master_clk_en;                                   // nios2_qsys_0:E_ci_multi_clk_en -> nios2_qsys_0_custom_instruction_master_translator:ci_slave_multi_clken
	wire   [4:0] nios2_qsys_0_custom_instruction_master_a;                                        // nios2_qsys_0:D_ci_a -> nios2_qsys_0_custom_instruction_master_translator:ci_slave_a
	wire   [7:0] nios2_qsys_0_custom_instruction_master_n;                                        // nios2_qsys_0:D_ci_n -> nios2_qsys_0_custom_instruction_master_translator:ci_slave_n
	wire         nios2_qsys_0_custom_instruction_master_writerc;                                  // nios2_qsys_0:D_ci_writerc -> nios2_qsys_0_custom_instruction_master_translator:ci_slave_writerc
	wire         nios2_qsys_0_custom_instruction_master_clk;                                      // nios2_qsys_0:E_ci_multi_clock -> nios2_qsys_0_custom_instruction_master_translator:ci_slave_multi_clk
	wire         nios2_qsys_0_custom_instruction_master_reset_req;                                // nios2_qsys_0:E_ci_multi_reset_req -> nios2_qsys_0_custom_instruction_master_translator:ci_slave_multi_reset_req
	wire         nios2_qsys_0_custom_instruction_master_start;                                    // nios2_qsys_0:E_ci_multi_start -> nios2_qsys_0_custom_instruction_master_translator:ci_slave_multi_start
	wire  [31:0] nios2_qsys_0_custom_instruction_master_dataa;                                    // nios2_qsys_0:E_ci_dataa -> nios2_qsys_0_custom_instruction_master_translator:ci_slave_dataa
	wire         nios2_qsys_0_custom_instruction_master_readra;                                   // nios2_qsys_0:D_ci_readra -> nios2_qsys_0_custom_instruction_master_translator:ci_slave_readra
	wire         nios2_qsys_0_custom_instruction_master_reset;                                    // nios2_qsys_0:E_ci_multi_reset -> nios2_qsys_0_custom_instruction_master_translator:ci_slave_multi_reset
	wire  [31:0] nios2_qsys_0_custom_instruction_master_datab;                                    // nios2_qsys_0:E_ci_datab -> nios2_qsys_0_custom_instruction_master_translator:ci_slave_datab
	wire         nios2_qsys_0_custom_instruction_master_readrb;                                   // nios2_qsys_0:D_ci_readrb -> nios2_qsys_0_custom_instruction_master_translator:ci_slave_readrb
	wire  [31:0] nios2_qsys_0_custom_instruction_master_translator_multi_ci_master_result;        // nios2_qsys_0_custom_instruction_master_multi_xconnect:ci_slave_result -> nios2_qsys_0_custom_instruction_master_translator:multi_ci_master_result
	wire   [4:0] nios2_qsys_0_custom_instruction_master_translator_multi_ci_master_b;             // nios2_qsys_0_custom_instruction_master_translator:multi_ci_master_b -> nios2_qsys_0_custom_instruction_master_multi_xconnect:ci_slave_b
	wire   [4:0] nios2_qsys_0_custom_instruction_master_translator_multi_ci_master_c;             // nios2_qsys_0_custom_instruction_master_translator:multi_ci_master_c -> nios2_qsys_0_custom_instruction_master_multi_xconnect:ci_slave_c
	wire   [4:0] nios2_qsys_0_custom_instruction_master_translator_multi_ci_master_a;             // nios2_qsys_0_custom_instruction_master_translator:multi_ci_master_a -> nios2_qsys_0_custom_instruction_master_multi_xconnect:ci_slave_a
	wire         nios2_qsys_0_custom_instruction_master_translator_multi_ci_master_clk_en;        // nios2_qsys_0_custom_instruction_master_translator:multi_ci_master_clken -> nios2_qsys_0_custom_instruction_master_multi_xconnect:ci_slave_clken
	wire         nios2_qsys_0_custom_instruction_master_translator_multi_ci_master_done;          // nios2_qsys_0_custom_instruction_master_multi_xconnect:ci_slave_done -> nios2_qsys_0_custom_instruction_master_translator:multi_ci_master_done
	wire   [7:0] nios2_qsys_0_custom_instruction_master_translator_multi_ci_master_n;             // nios2_qsys_0_custom_instruction_master_translator:multi_ci_master_n -> nios2_qsys_0_custom_instruction_master_multi_xconnect:ci_slave_n
	wire         nios2_qsys_0_custom_instruction_master_translator_multi_ci_master_writerc;       // nios2_qsys_0_custom_instruction_master_translator:multi_ci_master_writerc -> nios2_qsys_0_custom_instruction_master_multi_xconnect:ci_slave_writerc
	wire         nios2_qsys_0_custom_instruction_master_translator_multi_ci_master_clk;           // nios2_qsys_0_custom_instruction_master_translator:multi_ci_master_clk -> nios2_qsys_0_custom_instruction_master_multi_xconnect:ci_slave_clk
	wire         nios2_qsys_0_custom_instruction_master_translator_multi_ci_master_reset_req;     // nios2_qsys_0_custom_instruction_master_translator:multi_ci_master_reset_req -> nios2_qsys_0_custom_instruction_master_multi_xconnect:ci_slave_reset_req
	wire         nios2_qsys_0_custom_instruction_master_translator_multi_ci_master_start;         // nios2_qsys_0_custom_instruction_master_translator:multi_ci_master_start -> nios2_qsys_0_custom_instruction_master_multi_xconnect:ci_slave_start
	wire  [31:0] nios2_qsys_0_custom_instruction_master_translator_multi_ci_master_dataa;         // nios2_qsys_0_custom_instruction_master_translator:multi_ci_master_dataa -> nios2_qsys_0_custom_instruction_master_multi_xconnect:ci_slave_dataa
	wire         nios2_qsys_0_custom_instruction_master_translator_multi_ci_master_readra;        // nios2_qsys_0_custom_instruction_master_translator:multi_ci_master_readra -> nios2_qsys_0_custom_instruction_master_multi_xconnect:ci_slave_readra
	wire         nios2_qsys_0_custom_instruction_master_translator_multi_ci_master_reset;         // nios2_qsys_0_custom_instruction_master_translator:multi_ci_master_reset -> nios2_qsys_0_custom_instruction_master_multi_xconnect:ci_slave_reset
	wire  [31:0] nios2_qsys_0_custom_instruction_master_translator_multi_ci_master_datab;         // nios2_qsys_0_custom_instruction_master_translator:multi_ci_master_datab -> nios2_qsys_0_custom_instruction_master_multi_xconnect:ci_slave_datab
	wire         nios2_qsys_0_custom_instruction_master_translator_multi_ci_master_readrb;        // nios2_qsys_0_custom_instruction_master_translator:multi_ci_master_readrb -> nios2_qsys_0_custom_instruction_master_multi_xconnect:ci_slave_readrb
	wire  [31:0] nios2_qsys_0_custom_instruction_master_multi_xconnect_ci_master0_result;         // nios2_qsys_0_custom_instruction_master_multi_slave_translator0:ci_slave_result -> nios2_qsys_0_custom_instruction_master_multi_xconnect:ci_master0_result
	wire   [4:0] nios2_qsys_0_custom_instruction_master_multi_xconnect_ci_master0_b;              // nios2_qsys_0_custom_instruction_master_multi_xconnect:ci_master0_b -> nios2_qsys_0_custom_instruction_master_multi_slave_translator0:ci_slave_b
	wire   [4:0] nios2_qsys_0_custom_instruction_master_multi_xconnect_ci_master0_c;              // nios2_qsys_0_custom_instruction_master_multi_xconnect:ci_master0_c -> nios2_qsys_0_custom_instruction_master_multi_slave_translator0:ci_slave_c
	wire         nios2_qsys_0_custom_instruction_master_multi_xconnect_ci_master0_done;           // nios2_qsys_0_custom_instruction_master_multi_slave_translator0:ci_slave_done -> nios2_qsys_0_custom_instruction_master_multi_xconnect:ci_master0_done
	wire         nios2_qsys_0_custom_instruction_master_multi_xconnect_ci_master0_clk_en;         // nios2_qsys_0_custom_instruction_master_multi_xconnect:ci_master0_clken -> nios2_qsys_0_custom_instruction_master_multi_slave_translator0:ci_slave_clken
	wire   [4:0] nios2_qsys_0_custom_instruction_master_multi_xconnect_ci_master0_a;              // nios2_qsys_0_custom_instruction_master_multi_xconnect:ci_master0_a -> nios2_qsys_0_custom_instruction_master_multi_slave_translator0:ci_slave_a
	wire   [7:0] nios2_qsys_0_custom_instruction_master_multi_xconnect_ci_master0_n;              // nios2_qsys_0_custom_instruction_master_multi_xconnect:ci_master0_n -> nios2_qsys_0_custom_instruction_master_multi_slave_translator0:ci_slave_n
	wire         nios2_qsys_0_custom_instruction_master_multi_xconnect_ci_master0_writerc;        // nios2_qsys_0_custom_instruction_master_multi_xconnect:ci_master0_writerc -> nios2_qsys_0_custom_instruction_master_multi_slave_translator0:ci_slave_writerc
	wire  [31:0] nios2_qsys_0_custom_instruction_master_multi_xconnect_ci_master0_ipending;       // nios2_qsys_0_custom_instruction_master_multi_xconnect:ci_master0_ipending -> nios2_qsys_0_custom_instruction_master_multi_slave_translator0:ci_slave_ipending
	wire         nios2_qsys_0_custom_instruction_master_multi_xconnect_ci_master0_clk;            // nios2_qsys_0_custom_instruction_master_multi_xconnect:ci_master0_clk -> nios2_qsys_0_custom_instruction_master_multi_slave_translator0:ci_slave_clk
	wire         nios2_qsys_0_custom_instruction_master_multi_xconnect_ci_master0_reset_req;      // nios2_qsys_0_custom_instruction_master_multi_xconnect:ci_master0_reset_req -> nios2_qsys_0_custom_instruction_master_multi_slave_translator0:ci_slave_reset_req
	wire         nios2_qsys_0_custom_instruction_master_multi_xconnect_ci_master0_start;          // nios2_qsys_0_custom_instruction_master_multi_xconnect:ci_master0_start -> nios2_qsys_0_custom_instruction_master_multi_slave_translator0:ci_slave_start
	wire  [31:0] nios2_qsys_0_custom_instruction_master_multi_xconnect_ci_master0_dataa;          // nios2_qsys_0_custom_instruction_master_multi_xconnect:ci_master0_dataa -> nios2_qsys_0_custom_instruction_master_multi_slave_translator0:ci_slave_dataa
	wire         nios2_qsys_0_custom_instruction_master_multi_xconnect_ci_master0_readra;         // nios2_qsys_0_custom_instruction_master_multi_xconnect:ci_master0_readra -> nios2_qsys_0_custom_instruction_master_multi_slave_translator0:ci_slave_readra
	wire         nios2_qsys_0_custom_instruction_master_multi_xconnect_ci_master0_reset;          // nios2_qsys_0_custom_instruction_master_multi_xconnect:ci_master0_reset -> nios2_qsys_0_custom_instruction_master_multi_slave_translator0:ci_slave_reset
	wire  [31:0] nios2_qsys_0_custom_instruction_master_multi_xconnect_ci_master0_datab;          // nios2_qsys_0_custom_instruction_master_multi_xconnect:ci_master0_datab -> nios2_qsys_0_custom_instruction_master_multi_slave_translator0:ci_slave_datab
	wire         nios2_qsys_0_custom_instruction_master_multi_xconnect_ci_master0_readrb;         // nios2_qsys_0_custom_instruction_master_multi_xconnect:ci_master0_readrb -> nios2_qsys_0_custom_instruction_master_multi_slave_translator0:ci_slave_readrb
	wire         nios2_qsys_0_custom_instruction_master_multi_xconnect_ci_master0_estatus;        // nios2_qsys_0_custom_instruction_master_multi_xconnect:ci_master0_estatus -> nios2_qsys_0_custom_instruction_master_multi_slave_translator0:ci_slave_estatus
	wire  [31:0] nios2_qsys_0_custom_instruction_master_multi_slave_translator0_ci_master_result; // LCD_0:result -> nios2_qsys_0_custom_instruction_master_multi_slave_translator0:ci_master_result
	wire         nios2_qsys_0_custom_instruction_master_multi_slave_translator0_ci_master_start;  // nios2_qsys_0_custom_instruction_master_multi_slave_translator0:ci_master_start -> LCD_0:iniciar
	wire  [31:0] nios2_qsys_0_custom_instruction_master_multi_slave_translator0_ci_master_dataa;  // nios2_qsys_0_custom_instruction_master_multi_slave_translator0:ci_master_dataa -> LCD_0:dataA
	wire         nios2_qsys_0_custom_instruction_master_multi_slave_translator0_ci_master_done;   // LCD_0:done -> nios2_qsys_0_custom_instruction_master_multi_slave_translator0:ci_master_done
	wire         nios2_qsys_0_custom_instruction_master_multi_slave_translator0_ci_master_clk_en; // nios2_qsys_0_custom_instruction_master_multi_slave_translator0:ci_master_clken -> LCD_0:clk_en
	wire         nios2_qsys_0_custom_instruction_master_multi_slave_translator0_ci_master_reset;  // nios2_qsys_0_custom_instruction_master_multi_slave_translator0:ci_master_reset -> LCD_0:reset
	wire  [31:0] nios2_qsys_0_custom_instruction_master_multi_slave_translator0_ci_master_datab;  // nios2_qsys_0_custom_instruction_master_multi_slave_translator0:ci_master_datab -> LCD_0:dataB
	wire         nios2_qsys_0_custom_instruction_master_multi_slave_translator0_ci_master_clk;    // nios2_qsys_0_custom_instruction_master_multi_slave_translator0:ci_master_clk -> LCD_0:clk
	wire         nios2_qsys_0_data_master_waitrequest;                                            // mm_interconnect_0:nios2_qsys_0_data_master_waitrequest -> nios2_qsys_0:d_waitrequest
	wire  [31:0] nios2_qsys_0_data_master_writedata;                                              // nios2_qsys_0:d_writedata -> mm_interconnect_0:nios2_qsys_0_data_master_writedata
	wire  [13:0] nios2_qsys_0_data_master_address;                                                // nios2_qsys_0:d_address -> mm_interconnect_0:nios2_qsys_0_data_master_address
	wire         nios2_qsys_0_data_master_write;                                                  // nios2_qsys_0:d_write -> mm_interconnect_0:nios2_qsys_0_data_master_write
	wire         nios2_qsys_0_data_master_read;                                                   // nios2_qsys_0:d_read -> mm_interconnect_0:nios2_qsys_0_data_master_read
	wire  [31:0] nios2_qsys_0_data_master_readdata;                                               // mm_interconnect_0:nios2_qsys_0_data_master_readdata -> nios2_qsys_0:d_readdata
	wire         nios2_qsys_0_data_master_debugaccess;                                            // nios2_qsys_0:jtag_debug_module_debugaccess_to_roms -> mm_interconnect_0:nios2_qsys_0_data_master_debugaccess
	wire   [3:0] nios2_qsys_0_data_master_byteenable;                                             // nios2_qsys_0:d_byteenable -> mm_interconnect_0:nios2_qsys_0_data_master_byteenable
	wire         mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_waitrequest;                     // jtag_uart_0:av_waitrequest -> mm_interconnect_0:jtag_uart_0_avalon_jtag_slave_waitrequest
	wire  [31:0] mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_writedata;                       // mm_interconnect_0:jtag_uart_0_avalon_jtag_slave_writedata -> jtag_uart_0:av_writedata
	wire   [0:0] mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_address;                         // mm_interconnect_0:jtag_uart_0_avalon_jtag_slave_address -> jtag_uart_0:av_address
	wire         mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_chipselect;                      // mm_interconnect_0:jtag_uart_0_avalon_jtag_slave_chipselect -> jtag_uart_0:av_chipselect
	wire         mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_write;                           // mm_interconnect_0:jtag_uart_0_avalon_jtag_slave_write -> jtag_uart_0:av_write_n
	wire         mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_read;                            // mm_interconnect_0:jtag_uart_0_avalon_jtag_slave_read -> jtag_uart_0:av_read_n
	wire  [31:0] mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_readdata;                        // jtag_uart_0:av_readdata -> mm_interconnect_0:jtag_uart_0_avalon_jtag_slave_readdata
	wire         mm_interconnect_0_nios2_qsys_0_jtag_debug_module_waitrequest;                    // nios2_qsys_0:jtag_debug_module_waitrequest -> mm_interconnect_0:nios2_qsys_0_jtag_debug_module_waitrequest
	wire  [31:0] mm_interconnect_0_nios2_qsys_0_jtag_debug_module_writedata;                      // mm_interconnect_0:nios2_qsys_0_jtag_debug_module_writedata -> nios2_qsys_0:jtag_debug_module_writedata
	wire   [8:0] mm_interconnect_0_nios2_qsys_0_jtag_debug_module_address;                        // mm_interconnect_0:nios2_qsys_0_jtag_debug_module_address -> nios2_qsys_0:jtag_debug_module_address
	wire         mm_interconnect_0_nios2_qsys_0_jtag_debug_module_write;                          // mm_interconnect_0:nios2_qsys_0_jtag_debug_module_write -> nios2_qsys_0:jtag_debug_module_write
	wire         mm_interconnect_0_nios2_qsys_0_jtag_debug_module_read;                           // mm_interconnect_0:nios2_qsys_0_jtag_debug_module_read -> nios2_qsys_0:jtag_debug_module_read
	wire  [31:0] mm_interconnect_0_nios2_qsys_0_jtag_debug_module_readdata;                       // nios2_qsys_0:jtag_debug_module_readdata -> mm_interconnect_0:nios2_qsys_0_jtag_debug_module_readdata
	wire         mm_interconnect_0_nios2_qsys_0_jtag_debug_module_debugaccess;                    // mm_interconnect_0:nios2_qsys_0_jtag_debug_module_debugaccess -> nios2_qsys_0:jtag_debug_module_debugaccess
	wire   [3:0] mm_interconnect_0_nios2_qsys_0_jtag_debug_module_byteenable;                     // mm_interconnect_0:nios2_qsys_0_jtag_debug_module_byteenable -> nios2_qsys_0:jtag_debug_module_byteenable
	wire   [1:0] mm_interconnect_0_jumpbutton_s1_address;                                         // mm_interconnect_0:JumpButton_s1_address -> JumpButton:address
	wire  [31:0] mm_interconnect_0_jumpbutton_s1_readdata;                                        // JumpButton:readdata -> mm_interconnect_0:JumpButton_s1_readdata
	wire         nios2_qsys_0_instruction_master_waitrequest;                                     // mm_interconnect_0:nios2_qsys_0_instruction_master_waitrequest -> nios2_qsys_0:i_waitrequest
	wire  [13:0] nios2_qsys_0_instruction_master_address;                                         // nios2_qsys_0:i_address -> mm_interconnect_0:nios2_qsys_0_instruction_master_address
	wire         nios2_qsys_0_instruction_master_read;                                            // nios2_qsys_0:i_read -> mm_interconnect_0:nios2_qsys_0_instruction_master_read
	wire  [31:0] nios2_qsys_0_instruction_master_readdata;                                        // mm_interconnect_0:nios2_qsys_0_instruction_master_readdata -> nios2_qsys_0:i_readdata
	wire  [31:0] mm_interconnect_0_led_s1_writedata;                                              // mm_interconnect_0:LED_s1_writedata -> LED:writedata
	wire   [1:0] mm_interconnect_0_led_s1_address;                                                // mm_interconnect_0:LED_s1_address -> LED:address
	wire         mm_interconnect_0_led_s1_chipselect;                                             // mm_interconnect_0:LED_s1_chipselect -> LED:chipselect
	wire         mm_interconnect_0_led_s1_write;                                                  // mm_interconnect_0:LED_s1_write -> LED:write_n
	wire  [31:0] mm_interconnect_0_led_s1_readdata;                                               // LED:readdata -> mm_interconnect_0:LED_s1_readdata
	wire  [31:0] mm_interconnect_0_onchip_memory2_0_s1_writedata;                                 // mm_interconnect_0:onchip_memory2_0_s1_writedata -> onchip_memory2_0:writedata
	wire   [9:0] mm_interconnect_0_onchip_memory2_0_s1_address;                                   // mm_interconnect_0:onchip_memory2_0_s1_address -> onchip_memory2_0:address
	wire         mm_interconnect_0_onchip_memory2_0_s1_chipselect;                                // mm_interconnect_0:onchip_memory2_0_s1_chipselect -> onchip_memory2_0:chipselect
	wire         mm_interconnect_0_onchip_memory2_0_s1_clken;                                     // mm_interconnect_0:onchip_memory2_0_s1_clken -> onchip_memory2_0:clken
	wire         mm_interconnect_0_onchip_memory2_0_s1_write;                                     // mm_interconnect_0:onchip_memory2_0_s1_write -> onchip_memory2_0:write
	wire  [31:0] mm_interconnect_0_onchip_memory2_0_s1_readdata;                                  // onchip_memory2_0:readdata -> mm_interconnect_0:onchip_memory2_0_s1_readdata
	wire   [3:0] mm_interconnect_0_onchip_memory2_0_s1_byteenable;                                // mm_interconnect_0:onchip_memory2_0_s1_byteenable -> onchip_memory2_0:byteenable
	wire   [1:0] mm_interconnect_0_pausebutton_s1_address;                                        // mm_interconnect_0:PauseButton_s1_address -> PauseButton:address
	wire  [31:0] mm_interconnect_0_pausebutton_s1_readdata;                                       // PauseButton:readdata -> mm_interconnect_0:PauseButton_s1_readdata
	wire         irq_mapper_receiver0_irq;                                                        // jtag_uart_0:av_irq -> irq_mapper:receiver0_irq
	wire  [31:0] nios2_qsys_0_d_irq_irq;                                                          // irq_mapper:sender_irq -> nios2_qsys_0:d_irq
	wire         rst_controller_reset_out_reset;                                                  // rst_controller:reset_out -> [JumpButton:reset_n, LED:reset_n, PauseButton:reset_n, irq_mapper:reset, jtag_uart_0:rst_n, mm_interconnect_0:nios2_qsys_0_reset_n_reset_bridge_in_reset_reset, nios2_qsys_0:reset_n, onchip_memory2_0:reset, rst_translator:in_reset]
	wire         rst_controller_reset_out_reset_req;                                              // rst_controller:reset_req -> [nios2_qsys_0:reset_req, onchip_memory2_0:reset_req, rst_translator:reset_req_in]
	wire         nios2_qsys_0_jtag_debug_module_reset_reset;                                      // nios2_qsys_0:jtag_debug_module_resetrequest -> rst_controller:reset_in1

	CPU_nios2_qsys_0 nios2_qsys_0 (
		.clk                                   (clk_clk),                                                      //                       clk.clk
		.reset_n                               (~rst_controller_reset_out_reset),                              //                   reset_n.reset_n
		.reset_req                             (rst_controller_reset_out_reset_req),                           //                          .reset_req
		.d_address                             (nios2_qsys_0_data_master_address),                             //               data_master.address
		.d_byteenable                          (nios2_qsys_0_data_master_byteenable),                          //                          .byteenable
		.d_read                                (nios2_qsys_0_data_master_read),                                //                          .read
		.d_readdata                            (nios2_qsys_0_data_master_readdata),                            //                          .readdata
		.d_waitrequest                         (nios2_qsys_0_data_master_waitrequest),                         //                          .waitrequest
		.d_write                               (nios2_qsys_0_data_master_write),                               //                          .write
		.d_writedata                           (nios2_qsys_0_data_master_writedata),                           //                          .writedata
		.jtag_debug_module_debugaccess_to_roms (nios2_qsys_0_data_master_debugaccess),                         //                          .debugaccess
		.i_address                             (nios2_qsys_0_instruction_master_address),                      //        instruction_master.address
		.i_read                                (nios2_qsys_0_instruction_master_read),                         //                          .read
		.i_readdata                            (nios2_qsys_0_instruction_master_readdata),                     //                          .readdata
		.i_waitrequest                         (nios2_qsys_0_instruction_master_waitrequest),                  //                          .waitrequest
		.d_irq                                 (nios2_qsys_0_d_irq_irq),                                       //                     d_irq.irq
		.jtag_debug_module_resetrequest        (nios2_qsys_0_jtag_debug_module_reset_reset),                   //   jtag_debug_module_reset.reset
		.jtag_debug_module_address             (mm_interconnect_0_nios2_qsys_0_jtag_debug_module_address),     //         jtag_debug_module.address
		.jtag_debug_module_byteenable          (mm_interconnect_0_nios2_qsys_0_jtag_debug_module_byteenable),  //                          .byteenable
		.jtag_debug_module_debugaccess         (mm_interconnect_0_nios2_qsys_0_jtag_debug_module_debugaccess), //                          .debugaccess
		.jtag_debug_module_read                (mm_interconnect_0_nios2_qsys_0_jtag_debug_module_read),        //                          .read
		.jtag_debug_module_readdata            (mm_interconnect_0_nios2_qsys_0_jtag_debug_module_readdata),    //                          .readdata
		.jtag_debug_module_waitrequest         (mm_interconnect_0_nios2_qsys_0_jtag_debug_module_waitrequest), //                          .waitrequest
		.jtag_debug_module_write               (mm_interconnect_0_nios2_qsys_0_jtag_debug_module_write),       //                          .write
		.jtag_debug_module_writedata           (mm_interconnect_0_nios2_qsys_0_jtag_debug_module_writedata),   //                          .writedata
		.E_ci_multi_done                       (nios2_qsys_0_custom_instruction_master_done),                  // custom_instruction_master.done
		.E_ci_multi_clk_en                     (nios2_qsys_0_custom_instruction_master_clk_en),                //                          .clk_en
		.E_ci_multi_start                      (nios2_qsys_0_custom_instruction_master_start),                 //                          .start
		.E_ci_result                           (nios2_qsys_0_custom_instruction_master_result),                //                          .result
		.D_ci_a                                (nios2_qsys_0_custom_instruction_master_a),                     //                          .a
		.D_ci_b                                (nios2_qsys_0_custom_instruction_master_b),                     //                          .b
		.D_ci_c                                (nios2_qsys_0_custom_instruction_master_c),                     //                          .c
		.D_ci_n                                (nios2_qsys_0_custom_instruction_master_n),                     //                          .n
		.D_ci_readra                           (nios2_qsys_0_custom_instruction_master_readra),                //                          .readra
		.D_ci_readrb                           (nios2_qsys_0_custom_instruction_master_readrb),                //                          .readrb
		.D_ci_writerc                          (nios2_qsys_0_custom_instruction_master_writerc),               //                          .writerc
		.E_ci_dataa                            (nios2_qsys_0_custom_instruction_master_dataa),                 //                          .dataa
		.E_ci_datab                            (nios2_qsys_0_custom_instruction_master_datab),                 //                          .datab
		.E_ci_multi_clock                      (nios2_qsys_0_custom_instruction_master_clk),                   //                          .clk
		.E_ci_multi_reset                      (nios2_qsys_0_custom_instruction_master_reset),                 //                          .reset
		.E_ci_multi_reset_req                  (nios2_qsys_0_custom_instruction_master_reset_req)              //                          .reset_req
	);

	CPU_onchip_memory2_0 onchip_memory2_0 (
		.clk        (clk_clk),                                          //   clk1.clk
		.address    (mm_interconnect_0_onchip_memory2_0_s1_address),    //     s1.address
		.clken      (mm_interconnect_0_onchip_memory2_0_s1_clken),      //       .clken
		.chipselect (mm_interconnect_0_onchip_memory2_0_s1_chipselect), //       .chipselect
		.write      (mm_interconnect_0_onchip_memory2_0_s1_write),      //       .write
		.readdata   (mm_interconnect_0_onchip_memory2_0_s1_readdata),   //       .readdata
		.writedata  (mm_interconnect_0_onchip_memory2_0_s1_writedata),  //       .writedata
		.byteenable (mm_interconnect_0_onchip_memory2_0_s1_byteenable), //       .byteenable
		.reset      (rst_controller_reset_out_reset),                   // reset1.reset
		.reset_req  (rst_controller_reset_out_reset_req)                //       .reset_req
	);

	CPU_jtag_uart_0 jtag_uart_0 (
		.clk            (clk_clk),                                                     //               clk.clk
		.rst_n          (~rst_controller_reset_out_reset),                             //             reset.reset_n
		.av_chipselect  (mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_chipselect),  // avalon_jtag_slave.chipselect
		.av_address     (mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_address),     //                  .address
		.av_read_n      (~mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_read),       //                  .read_n
		.av_readdata    (mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_readdata),    //                  .readdata
		.av_write_n     (~mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_write),      //                  .write_n
		.av_writedata   (mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_writedata),   //                  .writedata
		.av_waitrequest (mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_waitrequest), //                  .waitrequest
		.av_irq         (irq_mapper_receiver0_irq)                                     //               irq.irq
	);

	display lcd_0 (
		.dataA   (nios2_qsys_0_custom_instruction_master_multi_slave_translator0_ci_master_dataa),  // nios_custom_instruction_slave.dataa
		.dataB   (nios2_qsys_0_custom_instruction_master_multi_slave_translator0_ci_master_datab),  //                              .datab
		.iniciar (nios2_qsys_0_custom_instruction_master_multi_slave_translator0_ci_master_start),  //                              .start
		.done    (nios2_qsys_0_custom_instruction_master_multi_slave_translator0_ci_master_done),   //                              .done
		.result  (nios2_qsys_0_custom_instruction_master_multi_slave_translator0_ci_master_result), //                              .result
		.clk_en  (nios2_qsys_0_custom_instruction_master_multi_slave_translator0_ci_master_clk_en), //                              .clk_en
		.clk     (nios2_qsys_0_custom_instruction_master_multi_slave_translator0_ci_master_clk),    //                              .clk
		.reset   (nios2_qsys_0_custom_instruction_master_multi_slave_translator0_ci_master_reset),  //                              .reset
		.rs      (lcd_0_conduit_end_export),                                                        //                   conduit_end.export
		.rw      (lcd_0_conduit_end_1_export),                                                      //                 conduit_end_1.export
		.enable  (lcd_0_conduit_end_2_export),                                                      //                 conduit_end_2.export
		.data    (lcd_0_conduit_end_3_export)                                                       //                 conduit_end_3.export
	);

	CPU_LED led (
		.clk        (clk_clk),                             //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),     //               reset.reset_n
		.address    (mm_interconnect_0_led_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_led_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_led_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_led_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_led_s1_readdata),   //                    .readdata
		.out_port   (led_external_connection_export)       // external_connection.export
	);

	CPU_JumpButton jumpbutton (
		.clk      (clk_clk),                                  //                 clk.clk
		.reset_n  (~rst_controller_reset_out_reset),          //               reset.reset_n
		.address  (mm_interconnect_0_jumpbutton_s1_address),  //                  s1.address
		.readdata (mm_interconnect_0_jumpbutton_s1_readdata), //                    .readdata
		.in_port  (jumpbutton_external_connection_export)     // external_connection.export
	);

	CPU_JumpButton pausebutton (
		.clk      (clk_clk),                                   //                 clk.clk
		.reset_n  (~rst_controller_reset_out_reset),           //               reset.reset_n
		.address  (mm_interconnect_0_pausebutton_s1_address),  //                  s1.address
		.readdata (mm_interconnect_0_pausebutton_s1_readdata), //                    .readdata
		.in_port  (pausebutton_external_connection_export)     // external_connection.export
	);

	altera_customins_master_translator #(
		.SHARED_COMB_AND_MULTI (1)
	) nios2_qsys_0_custom_instruction_master_translator (
		.ci_slave_dataa            (nios2_qsys_0_custom_instruction_master_dataa),                                //        ci_slave.dataa
		.ci_slave_datab            (nios2_qsys_0_custom_instruction_master_datab),                                //                .datab
		.ci_slave_result           (nios2_qsys_0_custom_instruction_master_result),                               //                .result
		.ci_slave_n                (nios2_qsys_0_custom_instruction_master_n),                                    //                .n
		.ci_slave_readra           (nios2_qsys_0_custom_instruction_master_readra),                               //                .readra
		.ci_slave_readrb           (nios2_qsys_0_custom_instruction_master_readrb),                               //                .readrb
		.ci_slave_writerc          (nios2_qsys_0_custom_instruction_master_writerc),                              //                .writerc
		.ci_slave_a                (nios2_qsys_0_custom_instruction_master_a),                                    //                .a
		.ci_slave_b                (nios2_qsys_0_custom_instruction_master_b),                                    //                .b
		.ci_slave_c                (nios2_qsys_0_custom_instruction_master_c),                                    //                .c
		.ci_slave_ipending         (),                                                                            //                .ipending
		.ci_slave_estatus          (),                                                                            //                .estatus
		.ci_slave_multi_clk        (nios2_qsys_0_custom_instruction_master_clk),                                  //                .clk
		.ci_slave_multi_reset      (nios2_qsys_0_custom_instruction_master_reset),                                //                .reset
		.ci_slave_multi_clken      (nios2_qsys_0_custom_instruction_master_clk_en),                               //                .clk_en
		.ci_slave_multi_reset_req  (nios2_qsys_0_custom_instruction_master_reset_req),                            //                .reset_req
		.ci_slave_multi_start      (nios2_qsys_0_custom_instruction_master_start),                                //                .start
		.ci_slave_multi_done       (nios2_qsys_0_custom_instruction_master_done),                                 //                .done
		.comb_ci_master_dataa      (),                                                                            //  comb_ci_master.dataa
		.comb_ci_master_datab      (),                                                                            //                .datab
		.comb_ci_master_result     (),                                                                            //                .result
		.comb_ci_master_n          (),                                                                            //                .n
		.comb_ci_master_readra     (),                                                                            //                .readra
		.comb_ci_master_readrb     (),                                                                            //                .readrb
		.comb_ci_master_writerc    (),                                                                            //                .writerc
		.comb_ci_master_a          (),                                                                            //                .a
		.comb_ci_master_b          (),                                                                            //                .b
		.comb_ci_master_c          (),                                                                            //                .c
		.comb_ci_master_ipending   (),                                                                            //                .ipending
		.comb_ci_master_estatus    (),                                                                            //                .estatus
		.multi_ci_master_clk       (nios2_qsys_0_custom_instruction_master_translator_multi_ci_master_clk),       // multi_ci_master.clk
		.multi_ci_master_reset     (nios2_qsys_0_custom_instruction_master_translator_multi_ci_master_reset),     //                .reset
		.multi_ci_master_clken     (nios2_qsys_0_custom_instruction_master_translator_multi_ci_master_clk_en),    //                .clk_en
		.multi_ci_master_reset_req (nios2_qsys_0_custom_instruction_master_translator_multi_ci_master_reset_req), //                .reset_req
		.multi_ci_master_start     (nios2_qsys_0_custom_instruction_master_translator_multi_ci_master_start),     //                .start
		.multi_ci_master_done      (nios2_qsys_0_custom_instruction_master_translator_multi_ci_master_done),      //                .done
		.multi_ci_master_dataa     (nios2_qsys_0_custom_instruction_master_translator_multi_ci_master_dataa),     //                .dataa
		.multi_ci_master_datab     (nios2_qsys_0_custom_instruction_master_translator_multi_ci_master_datab),     //                .datab
		.multi_ci_master_result    (nios2_qsys_0_custom_instruction_master_translator_multi_ci_master_result),    //                .result
		.multi_ci_master_n         (nios2_qsys_0_custom_instruction_master_translator_multi_ci_master_n),         //                .n
		.multi_ci_master_readra    (nios2_qsys_0_custom_instruction_master_translator_multi_ci_master_readra),    //                .readra
		.multi_ci_master_readrb    (nios2_qsys_0_custom_instruction_master_translator_multi_ci_master_readrb),    //                .readrb
		.multi_ci_master_writerc   (nios2_qsys_0_custom_instruction_master_translator_multi_ci_master_writerc),   //                .writerc
		.multi_ci_master_a         (nios2_qsys_0_custom_instruction_master_translator_multi_ci_master_a),         //                .a
		.multi_ci_master_b         (nios2_qsys_0_custom_instruction_master_translator_multi_ci_master_b),         //                .b
		.multi_ci_master_c         (nios2_qsys_0_custom_instruction_master_translator_multi_ci_master_c),         //                .c
		.ci_slave_multi_dataa      (32'b00000000000000000000000000000000),                                        //     (terminated)
		.ci_slave_multi_datab      (32'b00000000000000000000000000000000),                                        //     (terminated)
		.ci_slave_multi_result     (),                                                                            //     (terminated)
		.ci_slave_multi_n          (8'b00000000),                                                                 //     (terminated)
		.ci_slave_multi_readra     (1'b0),                                                                        //     (terminated)
		.ci_slave_multi_readrb     (1'b0),                                                                        //     (terminated)
		.ci_slave_multi_writerc    (1'b0),                                                                        //     (terminated)
		.ci_slave_multi_a          (5'b00000),                                                                    //     (terminated)
		.ci_slave_multi_b          (5'b00000),                                                                    //     (terminated)
		.ci_slave_multi_c          (5'b00000)                                                                     //     (terminated)
	);

	CPU_nios2_qsys_0_custom_instruction_master_multi_xconnect nios2_qsys_0_custom_instruction_master_multi_xconnect (
		.ci_slave_dataa       (nios2_qsys_0_custom_instruction_master_translator_multi_ci_master_dataa),     //   ci_slave.dataa
		.ci_slave_datab       (nios2_qsys_0_custom_instruction_master_translator_multi_ci_master_datab),     //           .datab
		.ci_slave_result      (nios2_qsys_0_custom_instruction_master_translator_multi_ci_master_result),    //           .result
		.ci_slave_n           (nios2_qsys_0_custom_instruction_master_translator_multi_ci_master_n),         //           .n
		.ci_slave_readra      (nios2_qsys_0_custom_instruction_master_translator_multi_ci_master_readra),    //           .readra
		.ci_slave_readrb      (nios2_qsys_0_custom_instruction_master_translator_multi_ci_master_readrb),    //           .readrb
		.ci_slave_writerc     (nios2_qsys_0_custom_instruction_master_translator_multi_ci_master_writerc),   //           .writerc
		.ci_slave_a           (nios2_qsys_0_custom_instruction_master_translator_multi_ci_master_a),         //           .a
		.ci_slave_b           (nios2_qsys_0_custom_instruction_master_translator_multi_ci_master_b),         //           .b
		.ci_slave_c           (nios2_qsys_0_custom_instruction_master_translator_multi_ci_master_c),         //           .c
		.ci_slave_ipending    (),                                                                            //           .ipending
		.ci_slave_estatus     (),                                                                            //           .estatus
		.ci_slave_clk         (nios2_qsys_0_custom_instruction_master_translator_multi_ci_master_clk),       //           .clk
		.ci_slave_reset       (nios2_qsys_0_custom_instruction_master_translator_multi_ci_master_reset),     //           .reset
		.ci_slave_clken       (nios2_qsys_0_custom_instruction_master_translator_multi_ci_master_clk_en),    //           .clk_en
		.ci_slave_reset_req   (nios2_qsys_0_custom_instruction_master_translator_multi_ci_master_reset_req), //           .reset_req
		.ci_slave_start       (nios2_qsys_0_custom_instruction_master_translator_multi_ci_master_start),     //           .start
		.ci_slave_done        (nios2_qsys_0_custom_instruction_master_translator_multi_ci_master_done),      //           .done
		.ci_master0_dataa     (nios2_qsys_0_custom_instruction_master_multi_xconnect_ci_master0_dataa),      // ci_master0.dataa
		.ci_master0_datab     (nios2_qsys_0_custom_instruction_master_multi_xconnect_ci_master0_datab),      //           .datab
		.ci_master0_result    (nios2_qsys_0_custom_instruction_master_multi_xconnect_ci_master0_result),     //           .result
		.ci_master0_n         (nios2_qsys_0_custom_instruction_master_multi_xconnect_ci_master0_n),          //           .n
		.ci_master0_readra    (nios2_qsys_0_custom_instruction_master_multi_xconnect_ci_master0_readra),     //           .readra
		.ci_master0_readrb    (nios2_qsys_0_custom_instruction_master_multi_xconnect_ci_master0_readrb),     //           .readrb
		.ci_master0_writerc   (nios2_qsys_0_custom_instruction_master_multi_xconnect_ci_master0_writerc),    //           .writerc
		.ci_master0_a         (nios2_qsys_0_custom_instruction_master_multi_xconnect_ci_master0_a),          //           .a
		.ci_master0_b         (nios2_qsys_0_custom_instruction_master_multi_xconnect_ci_master0_b),          //           .b
		.ci_master0_c         (nios2_qsys_0_custom_instruction_master_multi_xconnect_ci_master0_c),          //           .c
		.ci_master0_ipending  (nios2_qsys_0_custom_instruction_master_multi_xconnect_ci_master0_ipending),   //           .ipending
		.ci_master0_estatus   (nios2_qsys_0_custom_instruction_master_multi_xconnect_ci_master0_estatus),    //           .estatus
		.ci_master0_clk       (nios2_qsys_0_custom_instruction_master_multi_xconnect_ci_master0_clk),        //           .clk
		.ci_master0_reset     (nios2_qsys_0_custom_instruction_master_multi_xconnect_ci_master0_reset),      //           .reset
		.ci_master0_clken     (nios2_qsys_0_custom_instruction_master_multi_xconnect_ci_master0_clk_en),     //           .clk_en
		.ci_master0_reset_req (nios2_qsys_0_custom_instruction_master_multi_xconnect_ci_master0_reset_req),  //           .reset_req
		.ci_master0_start     (nios2_qsys_0_custom_instruction_master_multi_xconnect_ci_master0_start),      //           .start
		.ci_master0_done      (nios2_qsys_0_custom_instruction_master_multi_xconnect_ci_master0_done)        //           .done
	);

	altera_customins_slave_translator #(
		.N_WIDTH          (8),
		.USE_DONE         (1),
		.NUM_FIXED_CYCLES (0)
	) nios2_qsys_0_custom_instruction_master_multi_slave_translator0 (
		.ci_slave_dataa      (nios2_qsys_0_custom_instruction_master_multi_xconnect_ci_master0_dataa),          //  ci_slave.dataa
		.ci_slave_datab      (nios2_qsys_0_custom_instruction_master_multi_xconnect_ci_master0_datab),          //          .datab
		.ci_slave_result     (nios2_qsys_0_custom_instruction_master_multi_xconnect_ci_master0_result),         //          .result
		.ci_slave_n          (nios2_qsys_0_custom_instruction_master_multi_xconnect_ci_master0_n),              //          .n
		.ci_slave_readra     (nios2_qsys_0_custom_instruction_master_multi_xconnect_ci_master0_readra),         //          .readra
		.ci_slave_readrb     (nios2_qsys_0_custom_instruction_master_multi_xconnect_ci_master0_readrb),         //          .readrb
		.ci_slave_writerc    (nios2_qsys_0_custom_instruction_master_multi_xconnect_ci_master0_writerc),        //          .writerc
		.ci_slave_a          (nios2_qsys_0_custom_instruction_master_multi_xconnect_ci_master0_a),              //          .a
		.ci_slave_b          (nios2_qsys_0_custom_instruction_master_multi_xconnect_ci_master0_b),              //          .b
		.ci_slave_c          (nios2_qsys_0_custom_instruction_master_multi_xconnect_ci_master0_c),              //          .c
		.ci_slave_ipending   (nios2_qsys_0_custom_instruction_master_multi_xconnect_ci_master0_ipending),       //          .ipending
		.ci_slave_estatus    (nios2_qsys_0_custom_instruction_master_multi_xconnect_ci_master0_estatus),        //          .estatus
		.ci_slave_clk        (nios2_qsys_0_custom_instruction_master_multi_xconnect_ci_master0_clk),            //          .clk
		.ci_slave_clken      (nios2_qsys_0_custom_instruction_master_multi_xconnect_ci_master0_clk_en),         //          .clk_en
		.ci_slave_reset_req  (nios2_qsys_0_custom_instruction_master_multi_xconnect_ci_master0_reset_req),      //          .reset_req
		.ci_slave_reset      (nios2_qsys_0_custom_instruction_master_multi_xconnect_ci_master0_reset),          //          .reset
		.ci_slave_start      (nios2_qsys_0_custom_instruction_master_multi_xconnect_ci_master0_start),          //          .start
		.ci_slave_done       (nios2_qsys_0_custom_instruction_master_multi_xconnect_ci_master0_done),           //          .done
		.ci_master_dataa     (nios2_qsys_0_custom_instruction_master_multi_slave_translator0_ci_master_dataa),  // ci_master.dataa
		.ci_master_datab     (nios2_qsys_0_custom_instruction_master_multi_slave_translator0_ci_master_datab),  //          .datab
		.ci_master_result    (nios2_qsys_0_custom_instruction_master_multi_slave_translator0_ci_master_result), //          .result
		.ci_master_clk       (nios2_qsys_0_custom_instruction_master_multi_slave_translator0_ci_master_clk),    //          .clk
		.ci_master_clken     (nios2_qsys_0_custom_instruction_master_multi_slave_translator0_ci_master_clk_en), //          .clk_en
		.ci_master_reset     (nios2_qsys_0_custom_instruction_master_multi_slave_translator0_ci_master_reset),  //          .reset
		.ci_master_start     (nios2_qsys_0_custom_instruction_master_multi_slave_translator0_ci_master_start),  //          .start
		.ci_master_done      (nios2_qsys_0_custom_instruction_master_multi_slave_translator0_ci_master_done),   //          .done
		.ci_master_n         (),                                                                                // (terminated)
		.ci_master_readra    (),                                                                                // (terminated)
		.ci_master_readrb    (),                                                                                // (terminated)
		.ci_master_writerc   (),                                                                                // (terminated)
		.ci_master_a         (),                                                                                // (terminated)
		.ci_master_b         (),                                                                                // (terminated)
		.ci_master_c         (),                                                                                // (terminated)
		.ci_master_ipending  (),                                                                                // (terminated)
		.ci_master_estatus   (),                                                                                // (terminated)
		.ci_master_reset_req ()                                                                                 // (terminated)
	);

	CPU_mm_interconnect_0 mm_interconnect_0 (
		.clk_0_clk_clk                                    (clk_clk),                                                      //                                  clk_0_clk.clk
		.nios2_qsys_0_reset_n_reset_bridge_in_reset_reset (rst_controller_reset_out_reset),                               // nios2_qsys_0_reset_n_reset_bridge_in_reset.reset
		.nios2_qsys_0_data_master_address                 (nios2_qsys_0_data_master_address),                             //                   nios2_qsys_0_data_master.address
		.nios2_qsys_0_data_master_waitrequest             (nios2_qsys_0_data_master_waitrequest),                         //                                           .waitrequest
		.nios2_qsys_0_data_master_byteenable              (nios2_qsys_0_data_master_byteenable),                          //                                           .byteenable
		.nios2_qsys_0_data_master_read                    (nios2_qsys_0_data_master_read),                                //                                           .read
		.nios2_qsys_0_data_master_readdata                (nios2_qsys_0_data_master_readdata),                            //                                           .readdata
		.nios2_qsys_0_data_master_write                   (nios2_qsys_0_data_master_write),                               //                                           .write
		.nios2_qsys_0_data_master_writedata               (nios2_qsys_0_data_master_writedata),                           //                                           .writedata
		.nios2_qsys_0_data_master_debugaccess             (nios2_qsys_0_data_master_debugaccess),                         //                                           .debugaccess
		.nios2_qsys_0_instruction_master_address          (nios2_qsys_0_instruction_master_address),                      //            nios2_qsys_0_instruction_master.address
		.nios2_qsys_0_instruction_master_waitrequest      (nios2_qsys_0_instruction_master_waitrequest),                  //                                           .waitrequest
		.nios2_qsys_0_instruction_master_read             (nios2_qsys_0_instruction_master_read),                         //                                           .read
		.nios2_qsys_0_instruction_master_readdata         (nios2_qsys_0_instruction_master_readdata),                     //                                           .readdata
		.jtag_uart_0_avalon_jtag_slave_address            (mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_address),      //              jtag_uart_0_avalon_jtag_slave.address
		.jtag_uart_0_avalon_jtag_slave_write              (mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_write),        //                                           .write
		.jtag_uart_0_avalon_jtag_slave_read               (mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_read),         //                                           .read
		.jtag_uart_0_avalon_jtag_slave_readdata           (mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_readdata),     //                                           .readdata
		.jtag_uart_0_avalon_jtag_slave_writedata          (mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_writedata),    //                                           .writedata
		.jtag_uart_0_avalon_jtag_slave_waitrequest        (mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_waitrequest),  //                                           .waitrequest
		.jtag_uart_0_avalon_jtag_slave_chipselect         (mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_chipselect),   //                                           .chipselect
		.JumpButton_s1_address                            (mm_interconnect_0_jumpbutton_s1_address),                      //                              JumpButton_s1.address
		.JumpButton_s1_readdata                           (mm_interconnect_0_jumpbutton_s1_readdata),                     //                                           .readdata
		.LED_s1_address                                   (mm_interconnect_0_led_s1_address),                             //                                     LED_s1.address
		.LED_s1_write                                     (mm_interconnect_0_led_s1_write),                               //                                           .write
		.LED_s1_readdata                                  (mm_interconnect_0_led_s1_readdata),                            //                                           .readdata
		.LED_s1_writedata                                 (mm_interconnect_0_led_s1_writedata),                           //                                           .writedata
		.LED_s1_chipselect                                (mm_interconnect_0_led_s1_chipselect),                          //                                           .chipselect
		.nios2_qsys_0_jtag_debug_module_address           (mm_interconnect_0_nios2_qsys_0_jtag_debug_module_address),     //             nios2_qsys_0_jtag_debug_module.address
		.nios2_qsys_0_jtag_debug_module_write             (mm_interconnect_0_nios2_qsys_0_jtag_debug_module_write),       //                                           .write
		.nios2_qsys_0_jtag_debug_module_read              (mm_interconnect_0_nios2_qsys_0_jtag_debug_module_read),        //                                           .read
		.nios2_qsys_0_jtag_debug_module_readdata          (mm_interconnect_0_nios2_qsys_0_jtag_debug_module_readdata),    //                                           .readdata
		.nios2_qsys_0_jtag_debug_module_writedata         (mm_interconnect_0_nios2_qsys_0_jtag_debug_module_writedata),   //                                           .writedata
		.nios2_qsys_0_jtag_debug_module_byteenable        (mm_interconnect_0_nios2_qsys_0_jtag_debug_module_byteenable),  //                                           .byteenable
		.nios2_qsys_0_jtag_debug_module_waitrequest       (mm_interconnect_0_nios2_qsys_0_jtag_debug_module_waitrequest), //                                           .waitrequest
		.nios2_qsys_0_jtag_debug_module_debugaccess       (mm_interconnect_0_nios2_qsys_0_jtag_debug_module_debugaccess), //                                           .debugaccess
		.onchip_memory2_0_s1_address                      (mm_interconnect_0_onchip_memory2_0_s1_address),                //                        onchip_memory2_0_s1.address
		.onchip_memory2_0_s1_write                        (mm_interconnect_0_onchip_memory2_0_s1_write),                  //                                           .write
		.onchip_memory2_0_s1_readdata                     (mm_interconnect_0_onchip_memory2_0_s1_readdata),               //                                           .readdata
		.onchip_memory2_0_s1_writedata                    (mm_interconnect_0_onchip_memory2_0_s1_writedata),              //                                           .writedata
		.onchip_memory2_0_s1_byteenable                   (mm_interconnect_0_onchip_memory2_0_s1_byteenable),             //                                           .byteenable
		.onchip_memory2_0_s1_chipselect                   (mm_interconnect_0_onchip_memory2_0_s1_chipselect),             //                                           .chipselect
		.onchip_memory2_0_s1_clken                        (mm_interconnect_0_onchip_memory2_0_s1_clken),                  //                                           .clken
		.PauseButton_s1_address                           (mm_interconnect_0_pausebutton_s1_address),                     //                             PauseButton_s1.address
		.PauseButton_s1_readdata                          (mm_interconnect_0_pausebutton_s1_readdata)                     //                                           .readdata
	);

	CPU_irq_mapper irq_mapper (
		.clk           (clk_clk),                        //       clk.clk
		.reset         (rst_controller_reset_out_reset), // clk_reset.reset
		.receiver0_irq (irq_mapper_receiver0_irq),       // receiver0.irq
		.sender_irq    (nios2_qsys_0_d_irq_irq)          //    sender.irq
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (2),
		.OUTPUT_RESET_SYNC_EDGES   ("deassert"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (1),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller (
		.reset_in0      (~reset_reset_n),                             // reset_in0.reset
		.reset_in1      (nios2_qsys_0_jtag_debug_module_reset_reset), // reset_in1.reset
		.clk            (clk_clk),                                    //       clk.clk
		.reset_out      (rst_controller_reset_out_reset),             // reset_out.reset
		.reset_req      (rst_controller_reset_out_reset_req),         //          .reset_req
		.reset_req_in0  (1'b0),                                       // (terminated)
		.reset_req_in1  (1'b0),                                       // (terminated)
		.reset_in2      (1'b0),                                       // (terminated)
		.reset_req_in2  (1'b0),                                       // (terminated)
		.reset_in3      (1'b0),                                       // (terminated)
		.reset_req_in3  (1'b0),                                       // (terminated)
		.reset_in4      (1'b0),                                       // (terminated)
		.reset_req_in4  (1'b0),                                       // (terminated)
		.reset_in5      (1'b0),                                       // (terminated)
		.reset_req_in5  (1'b0),                                       // (terminated)
		.reset_in6      (1'b0),                                       // (terminated)
		.reset_req_in6  (1'b0),                                       // (terminated)
		.reset_in7      (1'b0),                                       // (terminated)
		.reset_req_in7  (1'b0),                                       // (terminated)
		.reset_in8      (1'b0),                                       // (terminated)
		.reset_req_in8  (1'b0),                                       // (terminated)
		.reset_in9      (1'b0),                                       // (terminated)
		.reset_req_in9  (1'b0),                                       // (terminated)
		.reset_in10     (1'b0),                                       // (terminated)
		.reset_req_in10 (1'b0),                                       // (terminated)
		.reset_in11     (1'b0),                                       // (terminated)
		.reset_req_in11 (1'b0),                                       // (terminated)
		.reset_in12     (1'b0),                                       // (terminated)
		.reset_req_in12 (1'b0),                                       // (terminated)
		.reset_in13     (1'b0),                                       // (terminated)
		.reset_req_in13 (1'b0),                                       // (terminated)
		.reset_in14     (1'b0),                                       // (terminated)
		.reset_req_in14 (1'b0),                                       // (terminated)
		.reset_in15     (1'b0),                                       // (terminated)
		.reset_req_in15 (1'b0)                                        // (terminated)
	);

endmodule
